
`timescale 1ns / 100ps

module widthReader(

   


   ) ;
   
   
   
   
endmodule